LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REGISTER_FILE IS
	PORT (
		OUT_REG_A : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		OUT_REG_B : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		INPUT_VAL : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		WRITE_ENABLE : IN STD_LOGIC;
		SEL_REG_A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEL_REG_B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		WRITE_REG_SEL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK : IN STD_LOGIC
	);
END REGISTER_FILE;

ARCHITECTURE Behavioral OF REGISTER_FILE IS
	TYPE REGISTER_FILE_TYPE IS ARRAY(0 TO 15) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL REGISTERS : REGISTER_FILE_TYPE;
BEGIN

	RegFile : PROCESS (CLK) IS
	BEGIN
		IF rising_edge(CLK) THEN
		
			-- Read A and B before bypass
			OUT_REG_A <= registers(to_integer(unsigned(SEL_REG_A)));
			OUT_REG_B <= registers(to_integer(unsigned(SEL_REG_B)));

			-- Write and bypass
			IF WRITE_ENABLE = '1' THEN
				registers(to_integer(unsigned(WRITE_REG_SEL))) <= INPUT_VAL; -- Write
				IF SEL_REG_A = WRITE_REG_SEL THEN -- Bypass for read A
          OUT_REG_A <= INPUT_VAL;
				END IF;
				IF SEL_REG_B = WRITE_REG_SEL THEN -- Bypass for read B
          OUT_REG_B <= INPUT_VAL;
				END IF;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;