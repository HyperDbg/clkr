LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TOP IS
	PORT (INPUT_CLK : IN STD_LOGIC_VECTOR (0 DOWNTO 0));
END TOP;

ARCHITECTURE Behavioral OF TOP IS

	-- RAM signals
	SIGNAL RAM_ADDR : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100"; 
	SIGNAL RAM_DATA_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM_WR : STD_LOGIC;
	SIGNAL RAM_CLOCK : STD_LOGIC; 
	SIGNAL RAM_DATA_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	-- RAM initialization signal
	SIGNAL IS_RAM_INITALIZED : STD_LOGIC := '0';
	SIGNAL PERFORM_RAM_INIT : STD_LOGIC := '0';

	-- Clock signal for testing purposes
	SIGNAL CLK : STD_LOGIC := '0';
	
	-- Instantiate components
	COMPONENT RAM
	PORT (
		RAM_ADDR : IN STD_LOGIC_VECTOR(6 DOWNTO 0); -- Address to write/read RAM
		RAM_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- Data to write into RAM
		RAM_WR : IN STD_LOGIC; -- Write enable
		RAM_CLOCK : IN STD_LOGIC; -- clock input for RAM
		RAM_DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) -- Data output of RAM
	);
	END COMPONENT;
	
	COMPONENT RAM_INIT 
	PORT (
		CLK : IN STD_LOGIC;
		PERFORM_INIT : IN STD_LOGIC
	);
	END COMPONENT;

BEGIN
	
	-- Using RAM
	RAM_UNT: RAM PORT MAP (RAM_ADDR => RAM_ADDR,
								  RAM_DATA_IN => RAM_DATA_IN,
								  RAM_WR => RAM_WR,
								  RAM_CLOCK => CLK,
								  RAM_DATA_OUT => RAM_DATA_OUT
								  );
								  
	-- Initialize RAM
	RAM_INITIALIZE: RAM_INIT PORT MAP (CLK => CLK,
								  PERFORM_INIT => PERFORM_RAM_INIT
								  );
								  
	PROCESS 
	BEGIN
		IF IS_RAM_INITALIZED = '0'
		THEN
			PERFORM_RAM_INIT <= '1';
		END IF;
	END PROCESS;
	
	-- Create testing signal
	PROCESS
	BEGIN
		CLK <= NOT CLK;
		WAIT FOR 1 ns;
	END PROCESS;

END Behavioral;